package tb_pkg;

    `include "wb_sim_master.sv"
    
endpackage