package tb_pkg;

    `include "wb_sim_master.sv"
    `include "mem/xpm_ram_model.sv"
    
endpackage